library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

-- Created from sslbp.bin
-- On 10/16/2013

entity sslbp is
	port (
	addra: in std_logic_vector(10 downto 0);
	addrb: in std_logic_vector(10 downto 0);
	clk: in std_logic;
	dina: in std_logic_vector(15 downto 0);
	douta: out std_logic_vector(15 downto 0);
	doutb: out std_logic_vector(15 downto 0);
	wea: in std_logic);
end sslbp;

architecture syn of sslbp is
   type ram_type is array (0 to 2047) of std_logic_vector(15 downto 0);
   signal RAM : ram_type := 
   (
   x"0000", x"0000", x"0000", x"0100", x"0800", x"0880", x"0100", x"B400",
   x"0C01", x"0480", x"0300", x"4006", x"B203", x"0101", x"B029", x"01FF",
   x"B02B", x"7234", x"B007", x"0138", x"B008", x"0149", x"B009", x"0132",
   x"B00A", x"0130", x"B00B", x"0137", x"B00C", x"0149", x"B00D", x"0136",
   x"B00E", x"0134", x"B00F", x"0112", x"B000", x"0101", x"B002", x"012B",
   x"B003", x"0108", x"B001", x"0170", x"B004", x"0132", x"B005", x"01D8",
   x"B006", x"0170", x"0800", x"0100", x"0880", x"0002", x"7007", x"B044",
   x"01A0", x"B42A", x"0125", x"B42B", x"0126", x"B42C", x"0100", x"B42D",
   x"0C32", x"0002", x"0002", x"01FF", x"C844", x"2038", x"0100", x"B04E",
   x"B200", x"7048", x"3617", x"704E", x"8052", x"8058", x"3616", x"7222",
   x"E05C", x"B065", x"7222", x"B05C", x"0170", x"0800", x"0100", x"0880",
   x"0180", x"0A00", x"0102", x"0A80", x"0100", x"0B00", x"0103", x"0B80",
   x"0101", x"B04F", x"01FE", x"B050", x"7007", x"B043", x"7052", x"A04F",
   x"308B", x"01FF", x"01C1", x"B413", x"66D9", x"0100", x"B410", x"B411",
   x"B412", x"B41D", x"B424", x"B720", x"B721", x"B723", x"B723", x"B740",
   x"B741", x"B742", x"B743", x"B760", x"B761", x"B762", x"B763", x"B640",
   x"B650", x"7050", x"A852", x"7050", x"A851", x"704F", x"8854", x"704F",
   x"8853", x"7050", x"A855", x"7051", x"A04F", x"35C4", x"0195", x"C410",
   x"0D80", x"0000", x"0000", x"0000", x"1800", x"11B2", x"11BB", x"11BF",
   x"11CB", x"11D1", x"1531", x"1539", x"11EC", x"11F4", x"11FB", x"1201",
   x"1209", x"121B", x"1221", x"1237", x"123D", x"1245", x"124D", x"1255",
   x"125D", x"1265", x"126D", x"1275", x"12AB", x"12DD", x"12E8", x"12F0",
   x"12FA", x"1301", x"1307", x"133B", x"134D", x"1358", x"1360", x"1367",
   x"136D", x"137A", x"1380", x"1388", x"139D", x"13AA", x"13B1", x"13BB",
   x"13C9", x"13D3", x"13DB", x"13ED", x"13FA", x"1401", x"140E", x"1415",
   x"141F", x"1427", x"1430", x"143A", x"1442", x"1455", x"1463", x"1117",
   x"112F", x"10D9", x"10EE", x"1173", x"1188", x"146A", x"14DE", x"1540",
   x"158D", x"7055", x"A04F", x"30ED", x"7411", x"8C12", x"0100", x"B411",
   x"6798", x"01BD", x"67B9", x"7720", x"67B9", x"7721", x"67B9", x"7722",
   x"67B9", x"7723", x"67BC", x"013D", x"B410", x"15C4", x"742E", x"6728",
   x"3110", x"7050", x"A855", x"7400", x"B740", x"7401", x"B741", x"7402",
   x"B742", x"7403", x"B743", x"8402", x"30FF", x"0101", x"8C13", x"7406",
   x"B720", x"7407", x"B721", x"7404", x"B722", x"7405", x"B723", x"7411",
   x"210B", x"7050", x"A856", x"7050", x"A857", x"013C", x"B410", x"1116",
   x"6775", x"5116", x"7050", x"A855", x"013C", x"B410", x"15C4", x"7411",
   x"8C12", x"0100", x"B411", x"704F", x"8858", x"6798", x"01BD", x"67B9",
   x"742F", x"B04D", x"312B", x"0003", x"0100", x"67B9", x"01FF", x"C84D",
   x"2124", x"0003", x"0003", x"67BE", x"013B", x"B410", x"15C4", x"742E",
   x"6728", x"3166", x"7222", x"E421", x"B430", x"017F", x"AC13", x"7050",
   x"A853", x"7050", x"A854", x"7055", x"A04F", x"3163", x"0114", x"C430",
   x"B423", x"0100", x"B400", x"B401", x"B402", x"B403", x"B404", x"B405",
   x"B406", x"B407", x"B408", x"B409", x"B40A", x"B40B", x"B40C", x"B40D",
   x"B40E", x"B40F", x"7424", x"3157", x"0142", x"B410", x"1162", x"0180",
   x"E41D", x"215D", x"013C", x"B410", x"1162", x"0174", x"E41D", x"2162",
   x"013E", x"B410", x"1165", x"013A", x"B410", x"1172", x"6775", x"5172",
   x"7055", x"A04F", x"316D", x"7050", x"A855", x"0180", x"A412", x"2172",
   x"013A", x"B410", x"15C4", x"7055", x"A04F", x"3187", x"7411", x"8C12",
   x"0100", x"B411", x"6798", x"01BD", x"67B9", x"7720", x"67B9", x"7721",
   x"67B9", x"7722", x"67B9", x"67B8", x"67BE", x"013F", x"B410", x"15C4",
   x"742E", x"6728", x"31AB", x"7050", x"A855", x"7400", x"B720", x"7401",
   x"B721", x"7402", x"B722", x"0108", x"A403", x"3198", x"0101", x"8C13",
   x"0100", x"B723", x"7404", x"B740", x"7405", x"B741", x"7406", x"B742",
   x"7407", x"B743", x"7411", x"21A6", x"7050", x"A856", x"7050", x"A857",
   x"013E", x"B410", x"11B1", x"6775", x"51B1", x"7050", x"A855", x"013E",
   x"B410", x"15C4", x"66D9", x"0100", x"B650", x"B640", x"0101", x"B410",
   x"7063", x"B423", x"15C4", x"67C3", x"0102", x"B410", x"15C4", x"7222",
   x"E421", x"B030", x"7223", x"F422", x"B031", x"7423", x"E030", x"41CA",
   x"0103", x"B410", x"15C4", x"6798", x"01DF", x"67BC", x"0104", x"B410",
   x"15C4", x"6775", x"51D6", x"0101", x"B410", x"11EB", x"0101", x"6728",
   x"31EB", x"015A", x"E400", x"21DF", x"0105", x"B410", x"11EB", x"7415",
   x"E41B", x"41E5", x"0101", x"CC15", x"11E7", x"0180", x"67E7", x"0102",
   x"67E7", x"0101", x"B410", x"15C4", x"6798", x"01E1", x"67B9", x"67B8",
   x"67BE", x"0108", x"B410", x"15C4", x"6727", x"31F9", x"0109", x"B410",
   x"11FA", x"6784", x"15C4", x"6798", x"01C1", x"67BC", x"010A", x"B410",
   x"15C4", x"0101", x"6728", x"3207", x"010B", x"B410", x"1208", x"6784",
   x"15C4", x"7400", x"220E", x"010C", x"B410", x"121A", x"0140", x"67E7",
   x"741A", x"E41B", x"4216", x"0101", x"CC1A", x"1218", x"0180", x"67E7",
   x"0101", x"B410", x"15C4", x"6798", x"01BC", x"67BC", x"010D", x"B410",
   x"15C4", x"0104", x"6728", x"322F", x"7400", x"B720", x"7401", x"B721",
   x"7402", x"B722", x"7403", x"B723", x"010E", x"B410", x"1236", x"6775",
   x"5236", x"010F", x"E047", x"2236", x"010E", x"B410", x"15C4", x"6798",
   x"01D0", x"67BC", x"010F", x"B410", x"15C4", x"0101", x"6728", x"3243",
   x"0110", x"B410", x"1244", x"6784", x"15C4", x"7400", x"B426", x"6798",
   x"01D1", x"67BC", x"0111", x"B410", x"15C4", x"0101", x"6728", x"3253",
   x"0112", x"B410", x"1254", x"6784", x"15C4", x"7400", x"B427", x"6798",
   x"01D2", x"67BC", x"0113", x"B410", x"15C4", x"0101", x"6728", x"3263",
   x"0114", x"B410", x"1264", x"6784", x"15C4", x"7400", x"B428", x"6798",
   x"01D3", x"67BC", x"0115", x"B410", x"15C4", x"0101", x"6728", x"3273",
   x"0116", x"B410", x"1274", x"6784", x"15C4", x"0117", x"B410", x"7426",
   x"B740", x"7427", x"B741", x"7428", x"B742", x"7400", x"B429", x"B743",
   x"7008", x"E426", x"B02F", x"0001", x"7009", x"F427", x"882F", x"0001",
   x"700A", x"F428", x"882F", x"0001", x"700B", x"F429", x"802F", x"22AA",
   x"0180", x"B41D", x"0108", x"B42E", x"0104", x"B42F", x"0109", x"E047",
   x"229D", x"01BF", x"AC13", x"0127", x"B410", x"010F", x"E047", x"22AA",
   x"013E", x"AC13", x"7050", x"A853", x"7050", x"A854", x"7064", x"B423",
   x"0140", x"B410", x"15C4", x"7400", x"B429", x"700C", x"E426", x"B02F",
   x"0001", x"700D", x"F427", x"882F", x"0001", x"700E", x"F428", x"882F",
   x"0001", x"700F", x"F429", x"802F", x"22D8", x"0174", x"B41D", x"0108",
   x"B42E", x"0104", x"B42F", x"0109", x"E047", x"22CA", x"01BE", x"AC13",
   x"0118", x"B410", x"010F", x"E047", x"22D7", x"013E", x"AC13", x"7050",
   x"A853", x"7050", x"A854", x"7064", x"B423", x"0140", x"B410", x"12DC",
   x"01FF", x"B424", x"011A", x"B410", x"15C4", x"6798", x"01BD", x"67B9",
   x"67B8", x"67B8", x"67B8", x"0108", x"67BC", x"0119", x"B410", x"15C4",
   x"742E", x"6728", x"32EE", x"013A", x"B410", x"12EF", x"6784", x"15C4",
   x"6798", x"01E6", x"67B9", x"7700", x"7703", x"67B9", x"67BE", x"011B",
   x"B410", x"15C4", x"6727", x"32FF", x"011C", x"B410", x"1300", x"6784",
   x"15C4", x"6798", x"01BB", x"67BC", x"011D", x"B410", x"15C4", x"0106",
   x"6728", x"332B", x"7400", x"B42E", x"7401", x"B42F", x"7402", x"B760",
   x"7403", x"B761", x"7404", x"B762", x"7405", x"B763", x"0109", x"E047",
   x"231D", x"01BF", x"AC13", x"011E", x"B410", x"010F", x"E047", x"232A",
   x"013E", x"AC13", x"7050", x"A853", x"7050", x"A854", x"7064", x"B423",
   x"0140", x"B410", x"133A", x"6775", x"533A", x"010F", x"E047", x"233A",
   x"013E", x"AC13", x"7050", x"A853", x"7050", x"A854", x"7064", x"B423",
   x"0140", x"B410", x"15C4", x"6798", x"01BD", x"67B9", x"742F", x"B04D",
   x"3349", x"0003", x"0100", x"67B9", x"01FF", x"C84D", x"2342", x"0003",
   x"0003", x"67BE", x"011F", x"B410", x"15C4", x"742E", x"6728", x"3353",
   x"0120", x"B410", x"1357", x"6775", x"5357", x"011E", x"B410", x"15C4",
   x"6798", x"01E7", x"67B9", x"67B6", x"67BE", x"0121", x"B410", x"15C4",
   x"6727", x"3365", x"0122", x"B410", x"1366", x"6784", x"15C4", x"6798",
   x"01C7", x"67BC", x"0123", x"B410", x"15C4", x"0101", x"6728", x"3378",
   x"7400", x"2375", x"0124", x"B410", x"1377", x"0122", x"B410", x"1379",
   x"6784", x"15C4", x"6798", x"01D7", x"67BC", x"0125", x"B410", x"15C4",
   x"0101", x"6728", x"3386", x"0126", x"B410", x"1387", x"6784", x"15C4",
   x"7400", x"238F", x"01FE", x"AC13", x"013A", x"B410", x"139C", x"B425",
   x"741A", x"E41B", x"4396", x"0101", x"CC1A", x"1398", x"0180", x"67E7",
   x"0140", x"67E7", x"0124", x"B410", x"15C4", x"6798", x"0165", x"67B9",
   x"0154", x"67B9", x"0108", x"67B9", x"67B6", x"67B6", x"67BE", x"0128",
   x"B410", x"15C4", x"6727", x"33AF", x"0129", x"B410", x"13B0", x"6784",
   x"15C4", x"6798", x"0145", x"67B9", x"0154", x"67B9", x"0108", x"67BC",
   x"012A", x"B410", x"15C4", x"0102", x"6728", x"33C7", x"7400", x"8401",
   x"23C4", x"012B", x"B410", x"13C6", x"0129", x"B410", x"13C8", x"6784",
   x"15C4", x"6798", x"0145", x"67B9", x"0152", x"67B9", x"0108", x"67BC",
   x"012C", x"B410", x"15C4", x"0102", x"6728", x"33D9", x"012D", x"B410",
   x"13DA", x"6784", x"15C4", x"7400", x"8401", x"B425", x"23E2", x"012E",
   x"B410", x"13EC", x"741A", x"E41B", x"43E8", x"0101", x"CC1A", x"13EA",
   x"0180", x"67E7", x"0140", x"67E7", x"15C4", x"6798", x"0165", x"67B9",
   x"0160", x"67B9", x"0108", x"67B9", x"67B8", x"67B8", x"67BE", x"012F",
   x"B410", x"15C4", x"6727", x"33FF", x"0130", x"B410", x"1400", x"6784",
   x"15C4", x"6798", x"0165", x"67B9", x"0104", x"67B9", x"0108", x"67B9",
   x"67B6", x"67B6", x"67BE", x"0131", x"B410", x"15C4", x"6727", x"3413",
   x"0132", x"B410", x"1414", x"6784", x"15C4", x"6798", x"0145", x"67B9",
   x"01FE", x"67B9", x"0108", x"67BC", x"0133", x"B410", x"15C4", x"0102",
   x"6728", x"3425", x"0134", x"B410", x"1426", x"6784", x"15C4", x"7400",
   x"8401", x"242D", x"0132", x"B410", x"142F", x"0135", x"B410", x"15C4",
   x"6798", x"0145", x"67B9", x"0152", x"67B9", x"0108", x"67BC", x"0136",
   x"B410", x"15C4", x"0102", x"6728", x"3440", x"0137", x"B410", x"1441",
   x"6784", x"15C4", x"7400", x"8401", x"244A", x"01FE", x"AC13", x"0138",
   x"B410", x"1454", x"741A", x"E41B", x"4450", x"0101", x"CC1A", x"1452",
   x"0180", x"67E7", x"0140", x"67E7", x"15C4", x"6798", x"0165", x"67B9",
   x"015C", x"67B9", x"0108", x"67B9", x"01F4", x"67B9", x"0101", x"67BC",
   x"0139", x"B410", x"15C4", x"6727", x"3468", x"013A", x"B410", x"1469",
   x"6784", x"15C4", x"7055", x"A04F", x"34DD", x"7411", x"8C12", x"0100",
   x"B411", x"7700", x"B04B", x"7703", x"B04A", x"7701", x"B04C", x"0140",
   x"A04A", x"247D", x"7050", x"A855", x"15C4", x"6798", x"704A", x"67B9",
   x"0103", x"A04A", x"B045", x"0001", x"0101", x"B046", x"7045", x"348D",
   x"01FF", x"C845", x"7046", x"C846", x"1486", x"01BF", x"E04A", x"54CF",
   x"0104", x"A04A", x"3498", x"0003", x"704B", x"67B9", x"704C", x"67B9",
   x"0120", x"A04A", x"34CC", x"0100", x"B41C", x"0108", x"E046", x"24B1",
   x"0003", x"7720", x"67B9", x"7721", x"67B9", x"7722", x"67B9", x"7723",
   x"67B9", x"7740", x"67B9", x"7741", x"67B9", x"7742", x"67B9", x"7743",
   x"67B9", x"0104", x"E046", x"24BD", x"0003", x"7720", x"67B9", x"7721",
   x"67B9", x"7722", x"67B9", x"7723", x"67B9", x"0102", x"E046", x"24C5",
   x"0003", x"7720", x"67B9", x"7721", x"67B9", x"0101", x"E046", x"24CB",
   x"0003", x"7720", x"67B9", x"14CE", x"7046", x"B41C", x"14DA", x"0120",
   x"A04A", x"34D8", x"0003", x"7720", x"67B9", x"0100", x"B41C", x"14DA",
   x"0101", x"B41C", x"67BE", x"0141", x"B410", x"15C4", x"741C", x"6728",
   x"352A", x"7050", x"A855", x"0108", x"E41C", x"24F6", x"7400", x"B720",
   x"7401", x"B721", x"7402", x"B722", x"7403", x"B723", x"7404", x"B740",
   x"7405", x"B741", x"7406", x"B742", x"7407", x"B743", x"0104", x"E41C",
   x"2506", x"7400", x"B720", x"7401", x"B721", x"7402", x"B722", x"7403",
   x"B723", x"0100", x"B740", x"B741", x"B742", x"B743", x"0102", x"E41C",
   x"2514", x"7400", x"B720", x"7401", x"B721", x"0100", x"B722", x"B723",
   x"B740", x"B741", x"B742", x"B743", x"0101", x"E41C", x"2521", x"7400",
   x"B720", x"0100", x"B721", x"B722", x"B723", x"B740", x"B741", x"B742",
   x"B743", x"7411", x"2525", x"7050", x"A856", x"7050", x"A857", x"0140",
   x"B410", x"1530", x"6775", x"5530", x"7050", x"A855", x"0140", x"B410",
   x"15C4", x"6798", x"01EB", x"67B9", x"0128", x"67BC", x"0106", x"B410",
   x"15C4", x"6727", x"353E", x"0107", x"B410", x"153F", x"6784", x"15C4",
   x"7055", x"A04F", x"358C", x"7411", x"8C12", x"0100", x"B411", x"742F",
   x"902B", x"0900", x"6798", x"01BD", x"67B9", x"742F", x"3589", x"0D02",
   x"7720", x"67B9", x"0500", x"3589", x"0D01", x"7721", x"67B9", x"0500",
   x"3589", x"0D01", x"7722", x"67B9", x"0500", x"3589", x"0D01", x"7723",
   x"67B9", x"0500", x"3589", x"0D01", x"7740", x"67B9", x"0500", x"3589",
   x"0D01", x"7741", x"67B9", x"0500", x"3589", x"0D01", x"7742", x"67B9",
   x"0500", x"3589", x"0D01", x"7743", x"67B9", x"0500", x"3589", x"0D01",
   x"7760", x"67B9", x"0500", x"3589", x"0D01", x"7761", x"67B9", x"0500",
   x"3589", x"0D01", x"7762", x"67B9", x"0500", x"3589", x"0003", x"7763",
   x"67B9", x"67BE", x"0143", x"B410", x"15C4", x"742E", x"6728", x"35BD",
   x"7050", x"A855", x"7400", x"B425", x"359A", x"0101", x"8C13", x"0140",
   x"67E7", x"159C", x"01BF", x"AC13", x"7401", x"B720", x"7402", x"B721",
   x"7403", x"B722", x"7404", x"B723", x"7405", x"B740", x"7406", x"B741",
   x"7407", x"B742", x"7408", x"B743", x"7409", x"B760", x"740A", x"B761",
   x"740B", x"B762", x"740C", x"B763", x"7411", x"25B8", x"7050", x"A856",
   x"7050", x"A857", x"0142", x"B410", x"15C3", x"6775", x"55C3", x"7050",
   x"A855", x"0142", x"B410", x"15C4", x"7412", x"B700", x"7413", x"B701",
   x"7410", x"B702", x"7425", x"B703", x"0C32", x"0E01", x"0F04", x"704F",
   x"C84F", x"902B", x"B050", x"01FF", x"C843", x"2066", x"0110", x"E04E",
   x"25EA", x"7053", x"902B", x"A051", x"A049", x"A055", x"A057", x"25EA",
   x"704F", x"8859", x"7050", x"A858", x"7056", x"B202", x"0100", x"B04E",
   x"B200", x"0001", x"0109", x"E04E", x"25FA", x"7054", x"A053", x"A049",
   x"25FA", x"7053", x"902B", x"A851", x"7053", x"B202", x"0100", x"B04E",
   x"B200", x"0001", x"010F", x"E04E", x"260A", x"7054", x"A053", x"A049",
   x"260A", x"7053", x"902B", x"A851", x"7053", x"B202", x"0100", x"B04E",
   x"B200", x"0001", x"0108", x"E04E", x"2616", x"7200", x"3616", x"7052",
   x"B202", x"A049", x"2616", x"0100", x"B04E", x"B200", x"166B", x"0100",
   x"B203", x"B047", x"01AA", x"B202", x"01FF", x"B052", x"0101", x"B04F",
   x"01FE", x"B050", x"0170", x"0800", x"0100", x"0880", x"0180", x"0A00",
   x"0102", x"0A80", x"0100", x"B049", x"7007", x"B044", x"01FF", x"C02B",
   x"7049", x"0200", x"B049", x"704F", x"C84F", x"902B", x"B050", x"742A",
   x"B034", x"742B", x"B035", x"742C", x"B036", x"742D", x"B037", x"66E4",
   x"66E4", x"66E4", x"66E4", x"0100", x"B032", x"B033", x"B038", x"B039",
   x"7230", x"B03A", x"7231", x"B03B", x"7232", x"B03C", x"7233", x"B03D",
   x"66ED", x"7032", x"B610", x"7033", x"B620", x"7034", x"B630", x"B640",
   x"0100", x"B650", x"0120", x"B670", x"0C32", x"0E01", x"01FF", x"C844",
   x"262E", x"01FF", x"B048", x"0108", x"E04E", x"266B", x"7200", x"266B",
   x"0100", x"B04E", x"B200", x"0101", x"A203", x"36D8", x"704E", x"26D2",
   x"7201", x"0980", x"B04E", x"7200", x"0900", x"B203", x"0110", x"A201",
   x"3682", x"7053", x"902B", x"A200", x"B055", x"B056", x"B057", x"01DE",
   x"AC13", x"16D1", x"0109", x"E201", x"269A", x"0120", x"B03A", x"01A1",
   x"B03B", x"0107", x"B03C", x"0100", x"B03D", x"67C8", x"01C8", x"B063",
   x"7201", x"B047", x"7051", x"902B", x"A200", x"B053", x"B054", x"7200",
   x"8851", x"16D1", x"0108", x"E201", x"26A3", x"7200", x"B052", x"26A2",
   x"0100", x"B048", x"16D1", x"010F", x"E201", x"26BD", x"0188", x"B03A",
   x"0113", x"B03B", x"0100", x"B03C", x"0100", x"B03D", x"67C8", x"0106",
   x"B063", x"01FA", x"B064", x"7201", x"B047", x"7051", x"902B", x"A200",
   x"B053", x"B054", x"7200", x"8851", x"16D1", x"0120", x"A201", x"36CC",
   x"0180", x"A201", x"36C6", x"7202", x"B580", x"16C8", x"7580", x"B202",
   x"0100", x"B04E", x"B200", x"16D1", x"01FF", x"B202", x"0100", x"B04E",
   x"B200", x"16D8", x"0108", x"E201", x"26D8", x"7201", x"B04E", x"B203",
   x"1049", x"0100", x"B414", x"B415", x"B416", x"B417", x"B418", x"B419",
   x"B41A", x"0114", x"B41B", x"1800", x"7034", x"C834", x"7035", x"D835",
   x"7036", x"D836", x"7037", x"D837", x"1800", x"0120", x"B03E", x"7032",
   x"C832", x"7033", x"D833", x"7034", x"D834", x"7035", x"D835", x"7036",
   x"D836", x"7037", x"D837", x"7038", x"D838", x"7039", x"D839", x"5719",
   x"7036", x"E03A", x"B036", x"7037", x"F03B", x"B037", x"7038", x"F03C",
   x"B038", x"7039", x"F03D", x"B039", x"4716", x"703A", x"C836", x"703B",
   x"D837", x"703C", x"D838", x"703D", x"D839", x"1718", x"0101", x"C832",
   x"1721", x"7036", x"E03A", x"B036", x"7037", x"F03B", x"B037", x"0101",
   x"C832", x"01FF", x"C83E", x"26EF", x"0003", x"0003", x"1800", x"0100",
   x"B02D", x"0D80", x"741E", x"2731", x"0C80", x"C029", x"B02E", x"B225",
   x"1738", x"0C80", x"3736", x"B02E", x"0001", x"1738", x"01FF", x"1800",
   x"7640", x"E02E", x"5773", x"0102", x"A650", x"374A", x"7419", x"E41B",
   x"4744", x"0101", x"CC19", x"1746", x"0180", x"67E7", x"0120", x"67E7",
   x"0100", x"1800", x"702D", x"375E", x"0400", x"B05A", x"0480", x"B05B",
   x"0003", x"0003", x"7600", x"B400", x"B224", x"0C01", x"01FF", x"C82D",
   x"2750", x"705A", x"0800", x"705B", x"0880", x"0003", x"741E", x"2770",
   x"7600", x"E224", x"376F", x"7414", x"E41B", x"4769", x"0101", x"CC14",
   x"176B", x"0180", x"67E7", x"0101", x"67E7", x"0100", x"1800", x"1771",
   x"C028", x"01FF", x"1774", x"0100", x"1800", x"7222", x"E421", x"E423",
   x"5800", x"7417", x"E41B", x"477F", x"0101", x"CC17", x"1781", x"0180",
   x"67E7", x"0108", x"67E7", x"1800", x"7222", x"E421", x"E423", x"5800",
   x"7417", x"E41B", x"478E", x"0101", x"CC17", x"1790", x"0180", x"67E7",
   x"0108", x"67E7", x"0180", x"A412", x"2797", x"0101", x"B410", x"1800",
   x"0003", x"7660", x"2798", x"B225", x"7640", x"37A8", x"7418", x"E41B",
   x"47A4", x"0101", x"CC18", x"17A6", x"0180", x"67E7", x"0110", x"67E7",
   x"0101", x"A640", x"37B5", x"7416", x"E41B", x"47B1", x"0101", x"CC16",
   x"17B3", x"0180", x"67E7", x"0104", x"67E7", x"1800", x"01FF", x"17B9",
   x"0100", x"B224", x"B600", x"1800", x"B224", x"B600", x"741E", x"27C3",
   x"0003", x"7224", x"B600", x"7222", x"B421", x"7223", x"B422", x"1800",
   x"7230", x"B032", x"7231", x"B033", x"7232", x"B034", x"7233", x"B035",
   x"0100", x"B036", x"B037", x"B038", x"B039", x"66ED", x"7032", x"B061",
   x"7033", x"B062", x"01FF", x"C861", x"01FF", x"D862", x"01FF", x"C861",
   x"01FF", x"D862", x"7061", x"B222", x"7062", x"B223", x"1800", x"8C12",
   x"7050", x"A857", x"0180", x"A412", x"37EF", x"7050", x"A854", x"0120",
   x"8C13", x"B640", x"0100", x"B650", x"1800", x"0000", x"0000", x"0000",
   x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"ABCD"
);

signal daddra: std_logic_vector(10 downto 0);
signal daddrb: std_logic_vector(10 downto 0);

begin
   asslbp: process (clk)
   begin
      if (clk'event and clk = '1') then
         if (wea = '1') then
            RAM(conv_integer(addra)) <= dina;
         end if;
         daddra <= addra;
         daddrb <= addrb;
      end if; -- clk 
   end process;

   douta <= RAM(conv_integer(daddra));
   doutb <= RAM(conv_integer(daddrb));
end;
